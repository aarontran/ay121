CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
240 130 30 200 9
0 70 1366 768
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 70 1366 768
144179218 0
0
6 Title:
5 Name:
0
0
0
15
10 Capacitor~
219 538 344 0 2 5
0 9 10
0
0 0 576 90
6 0.68�F
12 -5 54 3
2 Ce
14 -3 28 5
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
8953 0 0
0
0
9 Resistor~
219 510 344 0 3 5
0 2 12 -1
0
0 0 608 90
5 1.25k
7 -1 42 7
2 Rb
-20 -4 -6 4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4441 0 0
0
0
9 Resistor~
219 510 208 0 4 5
0 14 11 0 1
0
0 0 736 90
4 2.5k
6 -7 34 1
2 Rc
8 -6 22 2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3618 0 0
0
0
8 Speaker~
175 608 263 0 4 11
10 13 2 0 -1
0
0 0 4320 0
5 8 ohm
25 0 60 8
7 Speaker
19 -11 68 -3
0
0
11 %D %1 %2 %V
0
0
4 SIP2
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
3 SPK
6153 0 0
0
0
9 Resistor~
219 510 299 0 3 5
0 2 12 -1
0
0 0 608 90
5 1.25k
7 -1 42 7
2 Re
7 -3 21 5
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5394 0 0
0
0
9 Resistor~
219 465 226 0 4 5
0 10 4 0 1
0
0 0 96 90
3 22k
5 0 26 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7734 0 0
0
0
9 Resistor~
219 465 298 0 3 5
0 2 10 -1
0
0 0 224 90
3 13k
5 0 26 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9914 0 0
0
0
12 NPN Trans:C~
219 505 262 0 3 7
0 14 10 12
0
0 0 64 0
3 NPN
17 -3 38 5
2 Q1
21 -10 35 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
3747 0 0
0
0
10 Capacitor~
219 573 235 0 2 5
0 14 13
0
0 0 64 0
3 1�F
-9 -20 12 -12
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3549 0 0
0
0
7 Ground~
168 600 289 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7931 0 0
0
0
7 Ground~
168 510 380 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9325 0 0
0
0
2 +V
167 510 181 0 1 3
0 11
0
0 0 53600 0
3 +5V
-10 -14 11 -6
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8903 0 0
0
0
10 Capacitor~
219 438 262 0 2 5
0 9 10
0
0 0 64 0
6 0.68�F
-22 -20 20 -12
2 C2
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3834 0 0
0
0
7 Ground~
168 465 325 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3363 0 0
0
0
2 +V
167 465 199 0 1 3
0 4
0
0 0 53600 0
3 +5V
-10 -14 11 -6
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7668 0 0
0
0
15
1 0 0 0 0 0 0 11 0 0 2 2
510 374
510 362
1 1 0 0 0 0 0 1 2 0 0 3
538 353
538 362
510 362
1 2 0 0 0 0 0 5 2 0 0 2
510 317
510 326
2 2 0 0 0 0 0 1 2 0 0 3
538 335
538 326
510 326
1 2 4 0 0 0 0 15 6 0 0 2
465 208
465 208
1 1 2 0 0 0 0 14 7 0 0 4
465 319
465 321
465 321
465 316
2 0 10 0 0 0 0 7 0 0 8 2
465 280
465 262
1 0 10 0 0 0 0 6 0 0 9 2
465 244
465 262
2 2 10 0 0 0 0 13 8 0 0 2
447 262
487 262
1 2 11 0 0 0 0 12 3 0 0 2
510 190
510 190
2 3 12 0 0 0 0 5 8 0 0 4
510 281
510 284
510 284
510 280
1 2 2 0 0 0 0 10 4 0 0 2
600 283
600 279
1 2 13 0 0 0 0 4 9 0 0 3
600 247
600 235
582 235
1 0 14 0 0 0 0 9 0 0 15 2
564 235
510 235
1 1 14 0 0 0 0 3 8 0 0 2
510 226
510 244
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
