CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 100 30 200 9
0 70 1366 768
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 70 1366 768
8912914 32
0
6 Title:
5 Name:
0
0
0
27
2 +V
167 270 189 0 1 3
0 5
0
0 0 53600 0
3 +5V
-10 -14 11 -6
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8953 0 0
0
0
8 Antenna~
219 100 226 0 1 3
0 6
0
0 0 64 0
2 50
-8 -42 6 -34
4 ANT1
-14 -20 14 -12
0
0
10 %D %1 0 %V
0
0
3 BNC
3

0 1 1 0
82 0 0 0 1 0 0 0
3 ANT
4441 0 0
0
0
7 Ground~
168 270 315 0 1 3
0 2
0
0 0 53344 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3618 0 0
0
0
7 Ground~
168 176 306 0 1 3
0 2
0
0 0 53344 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6153 0 0
0
0
10 Capacitor~
219 243 252 0 2 5
0 3 7
0
0 0 320 180
3 1�F
-11 -20 10 -12
2 C5
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5394 0 0
0
0
10 Capacitor~
219 189 278 0 2 5
0 2 7
0
0 0 320 90
4 22nF
5 -14 33 -6
2 C4
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7734 0 0
0
0
7 Ground~
168 351 301 0 1 3
0 2
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9914 0 0
0
0
10 Capacitor~
219 351 279 0 2 5
0 2 9
0
0 0 320 90
5 100nF
-38 -14 -3 -6
2 C3
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3747 0 0
0
0
2 +V
167 432 189 0 1 3
0 4
0
0 0 53600 0
3 +5V
-10 -14 11 -6
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3549 0 0
0
0
7 Ground~
168 432 315 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7931 0 0
0
0
10 Capacitor~
219 405 252 0 2 5
0 9 10
0
0 0 320 0
6 0.68�F
-22 -20 20 -12
2 C2
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9325 0 0
0
0
2 +V
167 477 171 0 1 3
0 11
0
0 0 53600 0
3 +5V
-10 -14 11 -6
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8903 0 0
0
0
7 Ground~
168 477 315 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3834 0 0
0
0
7 Ground~
168 567 279 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3363 0 0
0
0
9 Inductor~
219 162 279 0 2 5
0 2 7
0
0 0 320 90
3 1�H
-32 -5 -11 3
2 L1
-28 -12 -14 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
7668 0 0
0
0
6 Diode~
219 288 252 0 2 5
0 3 8
0
0 0 64 0
5 DIODE
25 -51 60 -43
2 D1
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
4718 0 0
0
0
10 Capacitor~
219 540 225 0 2 5
0 14 13
0
0 0 320 0
3 1�F
-9 -20 12 -12
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3874 0 0
0
0
12 NPN Trans:C~
219 472 252 0 3 7
0 14 10 12
0
0 0 64 0
3 NPN
17 -3 38 5
2 Q1
21 -10 35 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
6671 0 0
0
0
9 Resistor~
219 144 252 0 2 5
0 7 6
0
0 0 352 180
2 33
-7 -14 7 -6
2 R8
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3789 0 0
0
0
9 Resistor~
219 270 288 0 4 5
0 3 2 0 -1
0
0 0 352 270
2 1k
8 -4 22 4
2 R7
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4871 0 0
0
0
9 Resistor~
219 270 219 0 3 5
0 5 3 1
0
0 0 352 270
4 6.3k
6 -3 34 5
2 R6
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3750 0 0
0
0
9 Resistor~
219 319 252 0 2 5
0 9 8
0
0 0 352 180
2 15
-7 -14 7 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8778 0 0
0
0
9 Resistor~
219 432 288 0 3 5
0 2 10 -1
0
0 0 352 90
3 13k
5 0 26 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
538 0 0
0
0
9 Resistor~
219 432 216 0 4 5
0 10 4 0 1
0
0 0 352 90
3 22k
5 0 26 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6843 0 0
0
0
9 Resistor~
219 477 289 0 3 5
0 2 12 -1
0
0 0 352 90
5 1.25k
7 -1 42 7
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3136 0 0
0
0
8 Speaker~
175 575 253 0 4 11
10 13 2 0 -1
0
0 0 4320 0
5 8 ohm
25 0 60 8
7 Speaker
19 -11 68 -3
0
0
11 %D %1 %2 %V
0
0
4 SIP2
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
3 SPK
5950 0 0
0
0
9 Resistor~
219 477 198 0 4 5
0 14 11 0 1
0
0 0 480 90
4 2.5k
6 -7 34 1
2 Re
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5670 0 0
0
0
27
1 0 3 0 0 4096 0 20 0 0 2 2
270 270
270 252
2 0 3 0 0 0 0 21 0 0 3 2
270 237
270 252
1 1 3 0 0 4224 0 5 16 0 0 2
252 252
278 252
1 2 4 0 0 0 0 9 24 0 0 2
432 198
432 198
1 1 5 0 0 4224 0 1 21 0 0 2
270 198
270 201
1 2 6 0 0 8320 0 2 19 0 0 3
100 242
100 252
126 252
1 0 2 0 0 4096 0 4 0 0 9 2
176 300
176 297
1 2 2 0 0 12288 0 3 20 0 0 4
270 309
270 311
270 311
270 306
1 1 2 0 0 4224 0 15 6 0 0 3
162 297
189 297
189 287
2 0 7 0 0 8192 0 6 0 0 11 3
189 269
189 261
176 261
0 2 7 0 0 8192 0 0 15 12 0 3
176 252
176 261
162 261
1 2 7 0 0 4224 0 19 5 0 0 2
162 252
234 252
2 2 8 0 0 4224 0 16 22 0 0 4
298 252
302 252
302 252
301 252
1 1 2 0 0 0 0 8 7 0 0 4
351 288
351 298
351 298
351 295
2 0 9 0 0 4096 0 8 0 0 16 2
351 270
351 252
1 1 9 0 0 4224 0 22 11 0 0 2
337 252
396 252
1 1 2 0 0 0 0 10 23 0 0 4
432 309
432 311
432 311
432 306
2 0 10 0 0 4096 0 23 0 0 19 2
432 270
432 252
1 0 10 0 0 0 0 24 0 0 20 2
432 234
432 252
2 2 10 0 0 4224 0 11 18 0 0 2
414 252
454 252
1 2 11 0 0 0 0 12 27 0 0 2
477 180
477 180
1 1 2 0 0 0 0 13 25 0 0 4
477 309
477 311
477 311
477 307
2 3 12 0 0 12416 0 25 18 0 0 4
477 271
477 274
477 274
477 270
1 2 2 0 0 0 0 14 26 0 0 2
567 273
567 269
1 2 13 0 0 8320 0 26 17 0 0 3
567 237
567 225
549 225
1 0 14 0 0 4224 0 17 0 0 27 2
531 225
477 225
1 1 14 0 0 0 0 27 18 0 0 2
477 216
477 234
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
